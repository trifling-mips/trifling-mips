`define REPL_TARGET 