`ifndef COMPILE_OPTIONS_SVH
`define COMPILE_OPTIONS_SVH

/**
	Options to control optional components to be compiled
	These options are used to speed up compilation when debugging
**/

// whether enable victim cache in write_buffer
`define VICTIM_CACHE_ENABLE

`endif
