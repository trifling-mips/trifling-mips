`ifndef INST_MM_SVH
`define INST_MM_SVH

/*
    This header defines common data structrue & constants in inst_mm module
*/

// cpu defs
`include "cpu_defs.svh"

`endif
