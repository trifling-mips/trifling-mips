// enable sim
`define REPL_SIM
