`ifndef REGS_SVH
`define REGS_SVH

/*
    This header defines common data structrue & constants in regs module
*/

// cpu defs
`include "cpu_defs.svh"

`endif
