`timescale 1us/1ns
`include "test_repl.svh"

module test_repl #(
	parameter int unsigned SET_ASSOC = 4
) (

);

