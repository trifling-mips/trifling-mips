`ifndef CPU_DEFS_SVH
`define CPU_DEFS_SVH

/*
	This header defines common data structrue & constants in cpu module
*/

// common defs
`include "cpu_defs.svh"

`endif
