`ifndef EXCEPT_SVH
`define EXCEPT_SVH

/*
    This header defines common data structrue & constants in except module
*/

// cpu defs
`include "cpu_defs.svh"

`endif
