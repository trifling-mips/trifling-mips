`ifndef CACHE_DEFS_SVH
`define CACHE_DEFS_SVH

/*
	This header defines common data structrue & constants in cache module
*/

// common defs
`include "common_defs.svh"

`endif
