`ifndef DECODE_SVH
`define DECODE_SVH

/*
    This header defines common data structrue & constants in decode module
*/

// cpu defs
`include "cpu_defs.svh"

`endif
