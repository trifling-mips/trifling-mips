`ifndef REPL_DEFS_SVH
`define REPL_DEFS_SVH

/*
    This header defines common data structrue & constants in repl module
*/

// cache defs
`include "cache_defs.svh"

// enable sim
// `define REPL_SIM

`endif
