`ifndef VICTIM_CACHE_SVH
`define VICTIM_CACHE_SVH

/*
    This header defines common data structrue & constants in victim_cache module
*/

// cache defs
`include "cache_defs.svh"

`endif
