`ifndef INST_DECODE_SVH
`define INST_DECODE_SVH

/*
    This header defines common data structrue & constants in inst_decode module
*/

// cpu defs
`include "cpu_defs.svh"

`endif
