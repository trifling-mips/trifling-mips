`ifndef CP0_SVH
`define CP0_SVH

/*
    This header defines common data structrue & constants in cp0 module
*/

// cpu defs
`include "cpu_defs.svh"

`endif
