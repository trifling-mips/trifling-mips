`ifndef TEST_CPU_SVH
`define TEST_CPU_SVH

/*
    This header defines common constants in test_cpu module
*/

// testbench_defs & cpu_defs
`include "testbench_defs.svh"
`include "cpu_defs.svh"

`endif
