`ifndef INST_EXEC_SVH
`define INST_EXEC_SVH

/*
    This header defines common data structrue & constants in inst_exec module
*/

// cpu defs
`include "cpu_defs.svh"

`endif
