`ifndef INST_FETCH_SVH
`define INST_FETCH_SVH

/*
    This header defines common data structrue & funs in inst_fetch module
*/

// cpu defs
`include "cpu_defs.svh"

`endif
